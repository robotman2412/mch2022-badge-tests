
module top (
    output wire my_ledinar
);
    
    assign my_ledinar = 1;
    
endmodule
